module sq_wave_gen (
    input clk,
    input next_sample,
    output [9:0] code
);
    assign code = 0;
endmodule
